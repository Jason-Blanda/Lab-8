module register(R,in,reset,clk);  
 output [31:0] R;  
 input [31:0] in;  
 input reset,clk;  
register reg0(R[0],in[0],reset,clk);  
 register reg1(R[1],in[1],reset,clk);  
 register reg2(R[2],in[2],reset,clk);  
 register reg3(R[3],in[3],reset,clk);  
 register reg4(R[4],in[4],reset,clk);  
 register reg5(R[5],in[5],reset,clk);  
 register reg6(R[6],in[6],reset,clk);  
 register reg7(R[7],in[7],reset,clk);  
 register reg8(R[8],in[8],reset,clk);  
 register reg9(R[9],in[9],reset,clk);  
 register reg10(R[10],in[10],reset,clk);  
 register reg11(R[11],in[11],reset,clk);  
 register reg12(R[12],in[12],reset,clk);  
 register reg13(R[13],in[13],reset,clk);  
 register reg14(R[14],in[14],reset,clk);  
 register reg15(R[15],in[15],reset,clk);  
 register reg16(R[16],in[16],reset,clk);  
 register reg17(R[17],in[17],reset,clk);  
 register reg18(R[18],in[18],reset,clk);  
 register reg19(R[19],in[19],reset,clk);  
 register reg20(R[20],in[20],reset,clk);  
 register reg21(R[21],in[21],reset,clk);  
 register reg22(R[22],in[22],reset,clk);  
 register reg23(R[23],in[23],reset,clk);  
 register reg24(R[24],in[24],reset,clk);  
 register reg25(R[25],in[25],reset,clk);  
 register reg26(R[26],in[26],reset,clk);  
 register reg27(R[27],in[27],reset,clk);  
 register reg28(R[28],in[28],reset,clk);  
 register reg29(R[29],in[29],reset,clk);  
 register reg30(R[30],in[30],reset,clk);  
 register reg31(R[31],in[31],reset,clk);  
 endmodule  
